module main

import os { input }

fn main() {
	name := input('Whats your name: ')
	println('Hello ' + name)
}
