module main

fn main() {
	mut msg := 'Hello World!'
	println(msg)

	msg = 'This is a new message'
	println(msg)
}
